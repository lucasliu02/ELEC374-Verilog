`timescale 1ns/10ps

module and_32_tb;
	reg  